module wave_display_tb(
	 
	 reg clk, reset;

    );


endmodule
